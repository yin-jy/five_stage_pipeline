
`include "DEFINE.v"
module InstructionMemory(
	input wire [`INST_ADDR_BUS] rom_addr_i,
	input wire rom_ce_i,
	output wire [`INST_BUS] rom_data_o
);
	
	assign rom_data_o=	(rom_ce_i==`CHIP_DISABLE)?`ZERO_WORD:
						(rom_addr_i==32'h00000000)?32'h08000003:
						(rom_addr_i==32'h00000004)?32'h080001af:
						(rom_addr_i==32'h00000008)?32'h080001c3:
						(rom_addr_i==32'h0000000C)?32'h3c01d091:
						(rom_addr_i==32'h00000010)?32'h3428bb44:
						(rom_addr_i==32'h00000014)?32'hac080000:
						(rom_addr_i==32'h00000018)?32'h3c01e7e1:
						(rom_addr_i==32'h0000001C)?32'h3429fafb:
						(rom_addr_i==32'h00000020)?32'hac090004:
						(rom_addr_i==32'h00000024)?32'h3c012082:
						(rom_addr_i==32'h00000028)?32'h342a353f:
						(rom_addr_i==32'h0000002C)?32'hac0a0008:
						(rom_addr_i==32'h00000030)?32'h3c01e9d3:
						(rom_addr_i==32'h00000034)?32'h342b0007:
						(rom_addr_i==32'h00000038)?32'hac0b000c:
						(rom_addr_i==32'h0000003C)?32'h3c01a1e2:
						(rom_addr_i==32'h00000040)?32'h342c4baa:
						(rom_addr_i==32'h00000044)?32'hac0c0010:
						(rom_addr_i==32'h00000048)?32'h3c0118f8:
						(rom_addr_i==32'h0000004C)?32'h342d6872:
						(rom_addr_i==32'h00000050)?32'hac0d0014:
						(rom_addr_i==32'h00000054)?32'h3c01474b:
						(rom_addr_i==32'h00000058)?32'h342ea8c6:
						(rom_addr_i==32'h0000005C)?32'hac0e0018:
						(rom_addr_i==32'h00000060)?32'h3c018c00:
						(rom_addr_i==32'h00000064)?32'h342f6d60:
						(rom_addr_i==32'h00000068)?32'hac0f001c:
						(rom_addr_i==32'h0000006C)?32'h3c01f51f:
						(rom_addr_i==32'h00000070)?32'h34282b00:
						(rom_addr_i==32'h00000074)?32'hac080020:
						(rom_addr_i==32'h00000078)?32'h3c01f702:
						(rom_addr_i==32'h0000007C)?32'h3429ef5f:
						(rom_addr_i==32'h00000080)?32'hac090024:
						(rom_addr_i==32'h00000084)?32'h3c012859:
						(rom_addr_i==32'h00000088)?32'h342a54b7:
						(rom_addr_i==32'h0000008C)?32'hac0a0028:
						(rom_addr_i==32'h00000090)?32'h3c01f878:
						(rom_addr_i==32'h00000094)?32'h342bc4bf:
						(rom_addr_i==32'h00000098)?32'hac0b002c:
						(rom_addr_i==32'h0000009C)?32'h3c01f508:
						(rom_addr_i==32'h000000A0)?32'h342ce4a4:
						(rom_addr_i==32'h000000A4)?32'hac0c0030:
						(rom_addr_i==32'h000000A8)?32'h3c017c41:
						(rom_addr_i==32'h000000AC)?32'h342d941a:
						(rom_addr_i==32'h000000B0)?32'hac0d0034:
						(rom_addr_i==32'h000000B4)?32'h3c01ccdf:
						(rom_addr_i==32'h000000B8)?32'h342e2e4a:
						(rom_addr_i==32'h000000BC)?32'hac0e0038:
						(rom_addr_i==32'h000000C0)?32'h3c012452:
						(rom_addr_i==32'h000000C4)?32'h342fa9c0:
						(rom_addr_i==32'h000000C8)?32'hac0f003c:
						(rom_addr_i==32'h000000CC)?32'h3c016bf8:
						(rom_addr_i==32'h000000D0)?32'h34288c24:
						(rom_addr_i==32'h000000D4)?32'hac080040:
						(rom_addr_i==32'h000000D8)?32'h3c01ea6d:
						(rom_addr_i==32'h000000DC)?32'h3429a4b4:
						(rom_addr_i==32'h000000E0)?32'hac090044:
						(rom_addr_i==32'h000000E4)?32'h3c01cace:
						(rom_addr_i==32'h000000E8)?32'h342a197c:
						(rom_addr_i==32'h000000EC)?32'hac0a0048:
						(rom_addr_i==32'h000000F0)?32'h3c01f5a1:
						(rom_addr_i==32'h000000F4)?32'h342b4bb0:
						(rom_addr_i==32'h000000F8)?32'hac0b004c:
						(rom_addr_i==32'h000000FC)?32'h3c01a7de:
						(rom_addr_i==32'h00000100)?32'h342c9f5a:
						(rom_addr_i==32'h00000104)?32'hac0c0050:
						(rom_addr_i==32'h00000108)?32'h3c010924:
						(rom_addr_i==32'h0000010C)?32'h342d668c:
						(rom_addr_i==32'h00000110)?32'hac0d0054:
						(rom_addr_i==32'h00000114)?32'h3c01d960:
						(rom_addr_i==32'h00000118)?32'h342e89c7:
						(rom_addr_i==32'h0000011C)?32'hac0e0058:
						(rom_addr_i==32'h00000120)?32'h3c01ef1a:
						(rom_addr_i==32'h00000124)?32'h342f2e76:
						(rom_addr_i==32'h00000128)?32'hac0f005c:
						(rom_addr_i==32'h0000012C)?32'h3c01adc1:
						(rom_addr_i==32'h00000130)?32'h3428964d:
						(rom_addr_i==32'h00000134)?32'hac080060:
						(rom_addr_i==32'h00000138)?32'h3c01c1fb:
						(rom_addr_i==32'h0000013C)?32'h342941d8:
						(rom_addr_i==32'h00000140)?32'hac090064:
						(rom_addr_i==32'h00000144)?32'h3c01be3d:
						(rom_addr_i==32'h00000148)?32'h342aedef:
						(rom_addr_i==32'h0000014C)?32'hac0a0068:
						(rom_addr_i==32'h00000150)?32'h3c016468:
						(rom_addr_i==32'h00000154)?32'h342bfd6e:
						(rom_addr_i==32'h00000158)?32'hac0b006c:
						(rom_addr_i==32'h0000015C)?32'h3c01a7cd:
						(rom_addr_i==32'h00000160)?32'h342c6626:
						(rom_addr_i==32'h00000164)?32'hac0c0070:
						(rom_addr_i==32'h00000168)?32'h3c012bd2:
						(rom_addr_i==32'h0000016C)?32'h342de40a:
						(rom_addr_i==32'h00000170)?32'hac0d0074:
						(rom_addr_i==32'h00000174)?32'h3c01b4bf:
						(rom_addr_i==32'h00000178)?32'h342e6fba:
						(rom_addr_i==32'h0000017C)?32'hac0e0078:
						(rom_addr_i==32'h00000180)?32'h3c010826:
						(rom_addr_i==32'h00000184)?32'h342f328a:
						(rom_addr_i==32'h00000188)?32'hac0f007c:
						(rom_addr_i==32'h0000018C)?32'h3c0146e4:
						(rom_addr_i==32'h00000190)?32'h34286cbc:
						(rom_addr_i==32'h00000194)?32'hac080080:
						(rom_addr_i==32'h00000198)?32'h3c010bd1:
						(rom_addr_i==32'h0000019C)?32'h3429e365:
						(rom_addr_i==32'h000001A0)?32'hac090084:
						(rom_addr_i==32'h000001A4)?32'h3c0118dd:
						(rom_addr_i==32'h000001A8)?32'h342aa0e0:
						(rom_addr_i==32'h000001AC)?32'hac0a0088:
						(rom_addr_i==32'h000001B0)?32'h3c01d2ce:
						(rom_addr_i==32'h000001B4)?32'h342b21da:
						(rom_addr_i==32'h000001B8)?32'hac0b008c:
						(rom_addr_i==32'h000001BC)?32'h3c01b1e0:
						(rom_addr_i==32'h000001C0)?32'h342c49e4:
						(rom_addr_i==32'h000001C4)?32'hac0c0090:
						(rom_addr_i==32'h000001C8)?32'h3c01512d:
						(rom_addr_i==32'h000001CC)?32'h342d6e78:
						(rom_addr_i==32'h000001D0)?32'hac0d0094:
						(rom_addr_i==32'h000001D4)?32'h3c01f341:
						(rom_addr_i==32'h000001D8)?32'h342ec090:
						(rom_addr_i==32'h000001DC)?32'hac0e0098:
						(rom_addr_i==32'h000001E0)?32'h3c0108d1:
						(rom_addr_i==32'h000001E4)?32'h342f7555:
						(rom_addr_i==32'h000001E8)?32'hac0f009c:
						(rom_addr_i==32'h000001EC)?32'h3c017051:
						(rom_addr_i==32'h000001F0)?32'h34288ce4:
						(rom_addr_i==32'h000001F4)?32'hac0800a0:
						(rom_addr_i==32'h000001F8)?32'h3c0161ad:
						(rom_addr_i==32'h000001FC)?32'h3429d0a7:
						(rom_addr_i==32'h00000200)?32'hac0900a4:
						(rom_addr_i==32'h00000204)?32'h3c01c3f8:
						(rom_addr_i==32'h00000208)?32'h342ae882:
						(rom_addr_i==32'h0000020C)?32'hac0a00a8:
						(rom_addr_i==32'h00000210)?32'h3c01cb92:
						(rom_addr_i==32'h00000214)?32'h342b3881:
						(rom_addr_i==32'h00000218)?32'hac0b00ac:
						(rom_addr_i==32'h0000021C)?32'h3c012fd6:
						(rom_addr_i==32'h00000220)?32'h342ce20d:
						(rom_addr_i==32'h00000224)?32'hac0c00b0:
						(rom_addr_i==32'h00000228)?32'h3c017d61:
						(rom_addr_i==32'h0000022C)?32'h342d330f:
						(rom_addr_i==32'h00000230)?32'hac0d00b4:
						(rom_addr_i==32'h00000234)?32'h3c017211:
						(rom_addr_i==32'h00000238)?32'h342eeff0:
						(rom_addr_i==32'h0000023C)?32'hac0e00b8:
						(rom_addr_i==32'h00000240)?32'h3c01a574:
						(rom_addr_i==32'h00000244)?32'h342fc4f9:
						(rom_addr_i==32'h00000248)?32'hac0f00bc:
						(rom_addr_i==32'h0000024C)?32'h3c01b598:
						(rom_addr_i==32'h00000250)?32'h3428eefd:
						(rom_addr_i==32'h00000254)?32'hac0800c0:
						(rom_addr_i==32'h00000258)?32'h3c01c133:
						(rom_addr_i==32'h0000025C)?32'h3429257a:
						(rom_addr_i==32'h00000260)?32'hac0900c4:
						(rom_addr_i==32'h00000264)?32'h3c0146a9:
						(rom_addr_i==32'h00000268)?32'h342a9457:
						(rom_addr_i==32'h0000026C)?32'hac0a00c8:
						(rom_addr_i==32'h00000270)?32'h3c01ae00:
						(rom_addr_i==32'h00000274)?32'h342bfea0:
						(rom_addr_i==32'h00000278)?32'hac0b00cc:
						(rom_addr_i==32'h0000027C)?32'h3c01a7b4:
						(rom_addr_i==32'h00000280)?32'h342c80b7:
						(rom_addr_i==32'h00000284)?32'hac0c00d0:
						(rom_addr_i==32'h00000288)?32'h3c0129a0:
						(rom_addr_i==32'h0000028C)?32'h342dec35:
						(rom_addr_i==32'h00000290)?32'hac0d00d4:
						(rom_addr_i==32'h00000294)?32'h3c011e76:
						(rom_addr_i==32'h00000298)?32'h342ea1cf:
						(rom_addr_i==32'h0000029C)?32'hac0e00d8:
						(rom_addr_i==32'h000002A0)?32'h3c017f94:
						(rom_addr_i==32'h000002A4)?32'h342fc959:
						(rom_addr_i==32'h000002A8)?32'hac0f00dc:
						(rom_addr_i==32'h000002AC)?32'h3c01f5b1:
						(rom_addr_i==32'h000002B0)?32'h3428c7b2:
						(rom_addr_i==32'h000002B4)?32'hac0800e0:
						(rom_addr_i==32'h000002B8)?32'h3c015723:
						(rom_addr_i==32'h000002BC)?32'h342984dc:
						(rom_addr_i==32'h000002C0)?32'hac0900e4:
						(rom_addr_i==32'h000002C4)?32'h3c0195d4:
						(rom_addr_i==32'h000002C8)?32'h342a1b7a:
						(rom_addr_i==32'h000002CC)?32'hac0a00e8:
						(rom_addr_i==32'h000002D0)?32'h3c01394b:
						(rom_addr_i==32'h000002D4)?32'h342bbd41:
						(rom_addr_i==32'h000002D8)?32'hac0b00ec:
						(rom_addr_i==32'h000002DC)?32'h3c01c053:
						(rom_addr_i==32'h000002E0)?32'h342c09ba:
						(rom_addr_i==32'h000002E4)?32'hac0c00f0:
						(rom_addr_i==32'h000002E8)?32'h3c01414d:
						(rom_addr_i==32'h000002EC)?32'h342de9da:
						(rom_addr_i==32'h000002F0)?32'hac0d00f4:
						(rom_addr_i==32'h000002F4)?32'h3c018186:
						(rom_addr_i==32'h000002F8)?32'h342e66be:
						(rom_addr_i==32'h000002FC)?32'hac0e00f8:
						(rom_addr_i==32'h00000300)?32'h3c01b2f6:
						(rom_addr_i==32'h00000304)?32'h342fb12d:
						(rom_addr_i==32'h00000308)?32'hac0f00fc:
						(rom_addr_i==32'h0000030C)?32'h3c01e412:
						(rom_addr_i==32'h00000310)?32'h34283c4e:
						(rom_addr_i==32'h00000314)?32'hac080100:
						(rom_addr_i==32'h00000318)?32'h3c01f594:
						(rom_addr_i==32'h0000031C)?32'h34291f73:
						(rom_addr_i==32'h00000320)?32'hac090104:
						(rom_addr_i==32'h00000324)?32'h3c018c16:
						(rom_addr_i==32'h00000328)?32'h342a5125:
						(rom_addr_i==32'h0000032C)?32'hac0a0108:
						(rom_addr_i==32'h00000330)?32'h3c01237c:
						(rom_addr_i==32'h00000334)?32'h342be438:
						(rom_addr_i==32'h00000338)?32'hac0b010c:
						(rom_addr_i==32'h0000033C)?32'h3c012638:
						(rom_addr_i==32'h00000340)?32'h342c21c7:
						(rom_addr_i==32'h00000344)?32'hac0c0110:
						(rom_addr_i==32'h00000348)?32'h3c0141ec:
						(rom_addr_i==32'h0000034C)?32'h342d0f9a:
						(rom_addr_i==32'h00000350)?32'hac0d0114:
						(rom_addr_i==32'h00000354)?32'h3c01d739:
						(rom_addr_i==32'h00000358)?32'h342e3f00:
						(rom_addr_i==32'h0000035C)?32'hac0e0118:
						(rom_addr_i==32'h00000360)?32'h3c014118:
						(rom_addr_i==32'h00000364)?32'h342fa30b:
						(rom_addr_i==32'h00000368)?32'hac0f011c:
						(rom_addr_i==32'h0000036C)?32'h3c01d074:
						(rom_addr_i==32'h00000370)?32'h3428f86a:
						(rom_addr_i==32'h00000374)?32'hac080120:
						(rom_addr_i==32'h00000378)?32'h3c013e57:
						(rom_addr_i==32'h0000037C)?32'h3429a700:
						(rom_addr_i==32'h00000380)?32'hac090124:
						(rom_addr_i==32'h00000384)?32'h3c01ede4:
						(rom_addr_i==32'h00000388)?32'h342a3887:
						(rom_addr_i==32'h0000038C)?32'hac0a0128:
						(rom_addr_i==32'h00000390)?32'h3c015998:
						(rom_addr_i==32'h00000394)?32'h342b893d:
						(rom_addr_i==32'h00000398)?32'hac0b012c:
						(rom_addr_i==32'h0000039C)?32'h3c013254:
						(rom_addr_i==32'h000003A0)?32'h342c10fb:
						(rom_addr_i==32'h000003A4)?32'hac0c0130:
						(rom_addr_i==32'h000003A8)?32'h3c014047:
						(rom_addr_i==32'h000003AC)?32'h342d081f:
						(rom_addr_i==32'h000003B0)?32'hac0d0134:
						(rom_addr_i==32'h000003B4)?32'h3c019db5:
						(rom_addr_i==32'h000003B8)?32'h342e1a99:
						(rom_addr_i==32'h000003BC)?32'hac0e0138:
						(rom_addr_i==32'h000003C0)?32'h3c017929:
						(rom_addr_i==32'h000003C4)?32'h342f7540:
						(rom_addr_i==32'h000003C8)?32'hac0f013c:
						(rom_addr_i==32'h000003CC)?32'h3c015a06:
						(rom_addr_i==32'h000003D0)?32'h34285b82:
						(rom_addr_i==32'h000003D4)?32'hac080140:
						(rom_addr_i==32'h000003D8)?32'h3c01d4b1:
						(rom_addr_i==32'h000003DC)?32'h34292f59:
						(rom_addr_i==32'h000003E0)?32'hac090144:
						(rom_addr_i==32'h000003E4)?32'h3c0195d3:
						(rom_addr_i==32'h000003E8)?32'h342ade13:
						(rom_addr_i==32'h000003EC)?32'hac0a0148:
						(rom_addr_i==32'h000003F0)?32'h3c018cba:
						(rom_addr_i==32'h000003F4)?32'h342bafb7:
						(rom_addr_i==32'h000003F8)?32'hac0b014c:
						(rom_addr_i==32'h000003FC)?32'h3c01eacd:
						(rom_addr_i==32'h00000400)?32'h342c3436:
						(rom_addr_i==32'h00000404)?32'hac0c0150:
						(rom_addr_i==32'h00000408)?32'h3c01492c:
						(rom_addr_i==32'h0000040C)?32'h342dbef6:
						(rom_addr_i==32'h00000410)?32'hac0d0154:
						(rom_addr_i==32'h00000414)?32'h3c01c1d7:
						(rom_addr_i==32'h00000418)?32'h342edfcd:
						(rom_addr_i==32'h0000041C)?32'hac0e0158:
						(rom_addr_i==32'h00000420)?32'h3c01c0f4:
						(rom_addr_i==32'h00000424)?32'h342f63d2:
						(rom_addr_i==32'h00000428)?32'hac0f015c:
						(rom_addr_i==32'h0000042C)?32'h3c016164:
						(rom_addr_i==32'h00000430)?32'h3428e627:
						(rom_addr_i==32'h00000434)?32'hac080160:
						(rom_addr_i==32'h00000438)?32'h3c01915c:
						(rom_addr_i==32'h0000043C)?32'h3429c251:
						(rom_addr_i==32'h00000440)?32'hac090164:
						(rom_addr_i==32'h00000444)?32'h3c01136b:
						(rom_addr_i==32'h00000448)?32'h342a2fcd:
						(rom_addr_i==32'h0000044C)?32'hac0a0168:
						(rom_addr_i==32'h00000450)?32'h3c010dcf:
						(rom_addr_i==32'h00000454)?32'h342baccb:
						(rom_addr_i==32'h00000458)?32'hac0b016c:
						(rom_addr_i==32'h0000045C)?32'h3c0187e2:
						(rom_addr_i==32'h00000460)?32'h342c5933:
						(rom_addr_i==32'h00000464)?32'hac0c0170:
						(rom_addr_i==32'h00000468)?32'h3c01c777:
						(rom_addr_i==32'h0000046C)?32'h342d80eb:
						(rom_addr_i==32'h00000470)?32'hac0d0174:
						(rom_addr_i==32'h00000474)?32'h3c01ef1b:
						(rom_addr_i==32'h00000478)?32'h342e52ff:
						(rom_addr_i==32'h0000047C)?32'hac0e0178:
						(rom_addr_i==32'h00000480)?32'h3c012141:
						(rom_addr_i==32'h00000484)?32'h342f8885:
						(rom_addr_i==32'h00000488)?32'hac0f017c:
						(rom_addr_i==32'h0000048C)?32'h3c01919e:
						(rom_addr_i==32'h00000490)?32'h34286d6d:
						(rom_addr_i==32'h00000494)?32'hac080180:
						(rom_addr_i==32'h00000498)?32'h3c017829:
						(rom_addr_i==32'h0000049C)?32'h3429fc2c:
						(rom_addr_i==32'h000004A0)?32'hac090184:
						(rom_addr_i==32'h000004A4)?32'h3c01030c:
						(rom_addr_i==32'h000004A8)?32'h342a0397:
						(rom_addr_i==32'h000004AC)?32'hac0a0188:
						(rom_addr_i==32'h000004B0)?32'h3c01564d:
						(rom_addr_i==32'h000004B4)?32'h342bab6c:
						(rom_addr_i==32'h000004B8)?32'hac0b018c:
						(rom_addr_i==32'h000004BC)?32'h3c012984:
						(rom_addr_i==32'h000004C0)?32'h342cc79e:
						(rom_addr_i==32'h000004C4)?32'hac0c0190:
						(rom_addr_i==32'h000004C8)?32'h3c01cb56:
						(rom_addr_i==32'h000004CC)?32'h342d3b4e:
						(rom_addr_i==32'h000004D0)?32'hac0d0194:
						(rom_addr_i==32'h000004D4)?32'h3c014fab:
						(rom_addr_i==32'h000004D8)?32'h342ec9fc:
						(rom_addr_i==32'h000004DC)?32'hac0e0198:
						(rom_addr_i==32'h000004E0)?32'h3c01874d:
						(rom_addr_i==32'h000004E4)?32'h342ff294:
						(rom_addr_i==32'h000004E8)?32'hac0f019c:
						(rom_addr_i==32'h000004EC)?32'h3c012a67:
						(rom_addr_i==32'h000004F0)?32'h3428f484:
						(rom_addr_i==32'h000004F4)?32'hac0801a0:
						(rom_addr_i==32'h000004F8)?32'h3c019a1b:
						(rom_addr_i==32'h000004FC)?32'h34297d0f:
						(rom_addr_i==32'h00000500)?32'hac0901a4:
						(rom_addr_i==32'h00000504)?32'h3c014352:
						(rom_addr_i==32'h00000508)?32'h342a160b:
						(rom_addr_i==32'h0000050C)?32'hac0a01a8:
						(rom_addr_i==32'h00000510)?32'h3c01a771:
						(rom_addr_i==32'h00000514)?32'h342bba51:
						(rom_addr_i==32'h00000518)?32'hac0b01ac:
						(rom_addr_i==32'h0000051C)?32'h3c01b070:
						(rom_addr_i==32'h00000520)?32'h342c5c97:
						(rom_addr_i==32'h00000524)?32'hac0c01b0:
						(rom_addr_i==32'h00000528)?32'h3c01bf86:
						(rom_addr_i==32'h0000052C)?32'h342ddce0:
						(rom_addr_i==32'h00000530)?32'hac0d01b4:
						(rom_addr_i==32'h00000534)?32'h3c017356:
						(rom_addr_i==32'h00000538)?32'h342eb1b7:
						(rom_addr_i==32'h0000053C)?32'hac0e01b8:
						(rom_addr_i==32'h00000540)?32'h3c011575:
						(rom_addr_i==32'h00000544)?32'h342f515d:
						(rom_addr_i==32'h00000548)?32'hac0f01bc:
						(rom_addr_i==32'h0000054C)?32'h3c013a9e:
						(rom_addr_i==32'h00000550)?32'h34283c10:
						(rom_addr_i==32'h00000554)?32'hac0801c0:
						(rom_addr_i==32'h00000558)?32'h3c01e9d0:
						(rom_addr_i==32'h0000055C)?32'h34297a32:
						(rom_addr_i==32'h00000560)?32'hac0901c4:
						(rom_addr_i==32'h00000564)?32'h3c012702:
						(rom_addr_i==32'h00000568)?32'h342a3ef0:
						(rom_addr_i==32'h0000056C)?32'hac0a01c8:
						(rom_addr_i==32'h00000570)?32'h3c01d368:
						(rom_addr_i==32'h00000574)?32'h342bbdcf:
						(rom_addr_i==32'h00000578)?32'hac0b01cc:
						(rom_addr_i==32'h0000057C)?32'h3c0189d0:
						(rom_addr_i==32'h00000580)?32'h342ccf51:
						(rom_addr_i==32'h00000584)?32'hac0c01d0:
						(rom_addr_i==32'h00000588)?32'h3c01ff02:
						(rom_addr_i==32'h0000058C)?32'h342daf4e:
						(rom_addr_i==32'h00000590)?32'hac0d01d4:
						(rom_addr_i==32'h00000594)?32'h3c011403:
						(rom_addr_i==32'h00000598)?32'h342e4fbb:
						(rom_addr_i==32'h0000059C)?32'hac0e01d8:
						(rom_addr_i==32'h000005A0)?32'h3c017153:
						(rom_addr_i==32'h000005A4)?32'h342f5cf3:
						(rom_addr_i==32'h000005A8)?32'hac0f01dc:
						(rom_addr_i==32'h000005AC)?32'h3c011b4d:
						(rom_addr_i==32'h000005B0)?32'h34289890:
						(rom_addr_i==32'h000005B4)?32'hac0801e0:
						(rom_addr_i==32'h000005B8)?32'h3c01f63e:
						(rom_addr_i==32'h000005BC)?32'h3429f3df:
						(rom_addr_i==32'h000005C0)?32'hac0901e4:
						(rom_addr_i==32'h000005C4)?32'h3c01012f:
						(rom_addr_i==32'h000005C8)?32'h342ab561:
						(rom_addr_i==32'h000005CC)?32'hac0a01e8:
						(rom_addr_i==32'h000005D0)?32'h3c01c660:
						(rom_addr_i==32'h000005D4)?32'h342b883f:
						(rom_addr_i==32'h000005D8)?32'hac0b01ec:
						(rom_addr_i==32'h000005DC)?32'h3c01d13a:
						(rom_addr_i==32'h000005E0)?32'h342cc8ac:
						(rom_addr_i==32'h000005E4)?32'hac0c01f0:
						(rom_addr_i==32'h000005E8)?32'h3c01de62:
						(rom_addr_i==32'h000005EC)?32'h342dc6b6:
						(rom_addr_i==32'h000005F0)?32'hac0d01f4:
						(rom_addr_i==32'h000005F4)?32'h3c01159d:
						(rom_addr_i==32'h000005F8)?32'h342e966b:
						(rom_addr_i==32'h000005FC)?32'hac0e01f8:
						(rom_addr_i==32'h00000600)?32'h3c016658:
						(rom_addr_i==32'h00000604)?32'h342f27db:
						(rom_addr_i==32'h00000608)?32'hac0f01fc:
						(rom_addr_i==32'h0000060C)?32'h3c014000:
						(rom_addr_i==32'h00000610)?32'h34280014:
						(rom_addr_i==32'h00000614)?32'h8d1b0000:
						(rom_addr_i==32'h00000618)?32'h20100080:
						(rom_addr_i==32'h0000061C)?32'h00008820:
						(rom_addr_i==32'h00000620)?32'h0230402a:
						(rom_addr_i==32'h00000624)?32'h1100000e:
						(rom_addr_i==32'h00000628)?32'h2632ffff:
						(rom_addr_i==32'h0000062C)?32'h0240402a:
						(rom_addr_i==32'h00000630)?32'h15000009:
						(rom_addr_i==32'h00000634)?32'h00124880:
						(rom_addr_i==32'h00000638)?32'h8d2a0000:
						(rom_addr_i==32'h0000063C)?32'h8d2b0004:
						(rom_addr_i==32'h00000640)?32'h016a402b:
						(rom_addr_i==32'h00000644)?32'h11000004:
						(rom_addr_i==32'h00000648)?32'had2a0004:
						(rom_addr_i==32'h0000064C)?32'had2b0000:
						(rom_addr_i==32'h00000650)?32'h2652ffff:
						(rom_addr_i==32'h00000654)?32'h0800018b:
						(rom_addr_i==32'h00000658)?32'h22310001:
						(rom_addr_i==32'h0000065C)?32'h08000188:
						(rom_addr_i==32'h00000660)?32'h3c014000:
						(rom_addr_i==32'h00000664)?32'h34280014:
						(rom_addr_i==32'h00000668)?32'h8d1e0000:
						(rom_addr_i==32'h0000066C)?32'h03dbd822:
						(rom_addr_i==32'h00000670)?32'h24100200:
						(rom_addr_i==32'h00000674)?32'h2408017f:
						(rom_addr_i==32'h00000678)?32'hae080000:
						(rom_addr_i==32'h0000067C)?32'h2409025b:
						(rom_addr_i==32'h00000680)?32'hae090004:
						(rom_addr_i==32'h00000684)?32'h240a046f:
						(rom_addr_i==32'h00000688)?32'hae0a0008:
						(rom_addr_i==32'h0000068C)?32'h240b084f:
						(rom_addr_i==32'h00000690)?32'hae0b000c:
						(rom_addr_i==32'h00000694)?32'h24110210:
						(rom_addr_i==32'h00000698)?32'hae3b0000:
						(rom_addr_i==32'h0000069C)?32'h3c014000:
						(rom_addr_i==32'h000006A0)?32'h34320010:
						(rom_addr_i==32'h000006A4)?32'h0c0001c4:
						(rom_addr_i==32'h000006A8)?32'h34191234:
						(rom_addr_i==32'h000006AC)?32'h34195678:
						(rom_addr_i==32'h000006B0)?32'h88888888://undefined instruction
						(rom_addr_i==32'h000006B4)?32'h080001ad:
						(rom_addr_i==32'h000006B8)?32'h00000000:
						(rom_addr_i==32'h000006BC)?32'h3c014000:
						(rom_addr_i==32'h000006C0)?32'h34280000:
						(rom_addr_i==32'h000006C4)?32'h8d090008:
						(rom_addr_i==32'h000006C8)?32'h3c01ffff:
						(rom_addr_i==32'h000006CC)?32'h3421fff9:
						(rom_addr_i==32'h000006D0)?32'h01214824:
						(rom_addr_i==32'h000006D4)?32'had090008:
						(rom_addr_i==32'h000006D8)?32'h0211402a:
						(rom_addr_i==32'h000006DC)?32'h11000002:
						(rom_addr_i==32'h000006E0)?32'h26100004:
						(rom_addr_i==32'h000006E4)?32'h080001bb:
						(rom_addr_i==32'h000006E8)?32'h2610fff4:
						(rom_addr_i==32'h000006EC)?32'h8e080000:
						(rom_addr_i==32'h000006F0)?32'hae480000:
						(rom_addr_i==32'h000006F4)?32'h3c014000:
						(rom_addr_i==32'h000006F8)?32'h34280000:
						(rom_addr_i==32'h000006FC)?32'h8d090008:
						(rom_addr_i==32'h00000700)?32'h35290002:
						(rom_addr_i==32'h00000704)?32'had090008:
						(rom_addr_i==32'h00000708)?32'h03400008:
						(rom_addr_i==32'h0000070C)?32'h080001c3:
						(rom_addr_i==32'h00000710)?32'h3c017fff:
						(rom_addr_i==32'h00000714)?32'h3421ffff:
						(rom_addr_i==32'h00000718)?32'h03e1f824:
						(rom_addr_i==32'h0000071C)?32'h3c014000:
						(rom_addr_i==32'h00000720)?32'h34280000:
						(rom_addr_i==32'h00000724)?32'had000008:
						(rom_addr_i==32'h00000728)?32'h2409d8ef:
						(rom_addr_i==32'h0000072C)?32'had090000:
						(rom_addr_i==32'h00000730)?32'had090004:
						(rom_addr_i==32'h00000734)?32'h20090003:
						(rom_addr_i==32'h00000738)?32'had090008:
						(rom_addr_i==32'h0000073C)?32'h03e00008:
						`ZERO_WORD;
endmodule
